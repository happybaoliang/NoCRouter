library verilog;
use verilog.vl_types.all;
entity tc_node_mac is
    generic(
        buffer_size     : integer := 32;
        num_message_classes: integer := 2;
        num_resource_classes: integer := 2;
        num_vcs_per_class: integer := 1;
        num_routers_per_dim: integer := 4;
        num_dimensions  : integer := 2;
        num_nodes_per_router: integer := 1;
        connectivity    : integer := 0;
        packet_format   : integer := 2;
        flow_ctrl_type  : integer := 0;
        flow_ctrl_bypass: integer := 1;
        max_payload_length: integer := 4;
        min_payload_length: integer := 1;
        enable_link_pm  : integer := 1;
        flit_data_width : integer := 64;
        error_capture_mode: integer := 1;
        routing_type    : integer := 0;
        dim_order       : integer := 0;
        fb_mgmt_type    : integer := 0;
        disable_static_reservations: integer := 0;
        elig_mask       : integer := 0;
        lfsr_index      : integer := 0;
        cfg_node_addr_width: integer := 10;
        cfg_reg_addr_width: integer := 6;
        num_cfg_node_addrs: integer := 2;
        cfg_data_width  : integer := 32;
        num_packets_width: integer := 20;
        arrival_rv_width: integer := 20;
        mc_idx_rv_width : integer := 1;
        rc_idx_rv_width : integer := 1;
        plength_idx_rv_width: integer := 1;
        num_plength_vals: integer := 2;
        packet_count_width: integer := 8;
        reset_type      : integer := 0
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        address         : in     vl_logic_vector;
        channel_out     : out    vl_logic_vector;
        flow_ctrl_in    : in     vl_logic_vector;
        channel_in      : in     vl_logic_vector;
        flow_ctrl_out   : out    vl_logic_vector;
        cfg_node_addrs  : in     vl_logic_vector;
        cfg_req         : in     vl_logic;
        cfg_write       : in     vl_logic;
        cfg_addr        : in     vl_logic_vector;
        cfg_write_data  : in     vl_logic_vector;
        cfg_read_data   : out    vl_logic_vector;
        cfg_done        : out    vl_logic;
        error           : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of buffer_size : constant is 1;
    attribute mti_svvh_generic_type of num_message_classes : constant is 1;
    attribute mti_svvh_generic_type of num_resource_classes : constant is 1;
    attribute mti_svvh_generic_type of num_vcs_per_class : constant is 1;
    attribute mti_svvh_generic_type of num_routers_per_dim : constant is 1;
    attribute mti_svvh_generic_type of num_dimensions : constant is 1;
    attribute mti_svvh_generic_type of num_nodes_per_router : constant is 1;
    attribute mti_svvh_generic_type of connectivity : constant is 1;
    attribute mti_svvh_generic_type of packet_format : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_type : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_bypass : constant is 1;
    attribute mti_svvh_generic_type of max_payload_length : constant is 1;
    attribute mti_svvh_generic_type of min_payload_length : constant is 1;
    attribute mti_svvh_generic_type of enable_link_pm : constant is 1;
    attribute mti_svvh_generic_type of flit_data_width : constant is 1;
    attribute mti_svvh_generic_type of error_capture_mode : constant is 1;
    attribute mti_svvh_generic_type of routing_type : constant is 1;
    attribute mti_svvh_generic_type of dim_order : constant is 1;
    attribute mti_svvh_generic_type of fb_mgmt_type : constant is 1;
    attribute mti_svvh_generic_type of disable_static_reservations : constant is 1;
    attribute mti_svvh_generic_type of elig_mask : constant is 1;
    attribute mti_svvh_generic_type of lfsr_index : constant is 1;
    attribute mti_svvh_generic_type of cfg_node_addr_width : constant is 1;
    attribute mti_svvh_generic_type of cfg_reg_addr_width : constant is 1;
    attribute mti_svvh_generic_type of num_cfg_node_addrs : constant is 1;
    attribute mti_svvh_generic_type of cfg_data_width : constant is 1;
    attribute mti_svvh_generic_type of num_packets_width : constant is 1;
    attribute mti_svvh_generic_type of arrival_rv_width : constant is 1;
    attribute mti_svvh_generic_type of mc_idx_rv_width : constant is 1;
    attribute mti_svvh_generic_type of rc_idx_rv_width : constant is 1;
    attribute mti_svvh_generic_type of plength_idx_rv_width : constant is 1;
    attribute mti_svvh_generic_type of num_plength_vals : constant is 1;
    attribute mti_svvh_generic_type of packet_count_width : constant is 1;
    attribute mti_svvh_generic_type of reset_type : constant is 1;
end tc_node_mac;
