library verilog;
use verilog.vl_types.all;
entity tc_router_wrap is
    generic(
        topology        : integer := 0;
        buffer_size     : integer := 16;
        num_message_classes: integer := 2;
        num_resource_classes: integer := 1;
        num_vcs_per_class: integer := 1;
        num_nodes       : integer := 64;
        num_dimensions  : integer := 2;
        num_nodes_per_router: integer := 1;
        packet_format   : integer := 2;
        flow_ctrl_type  : integer := 0;
        flow_ctrl_bypass: integer := 0;
        max_payload_length: integer := 4;
        min_payload_length: integer := 0;
        router_type     : integer := 1;
        enable_link_pm  : integer := 1;
        flit_data_width : integer := 64;
        error_capture_mode: integer := 1;
        restrict_turns  : integer := 1;
        predecode_lar_info: integer := 1;
        routing_type    : integer := 0;
        dim_order       : integer := 0;
        input_stage_can_hold: integer := 0;
        fb_regfile_type : integer := 0;
        fb_mgmt_type    : integer := 0;
        fb_fast_peek    : integer := 1;
        disable_static_reservations: integer := 0;
        explicit_pipeline_register: integer := 1;
        gate_buffer_write: integer := 0;
        dual_path_alloc : integer := 0;
        dual_path_allow_conflicts: integer := 0;
        dual_path_mask_on_ready: integer := 1;
        precomp_ivc_sel : integer := 0;
        precomp_ip_sel  : integer := 0;
        elig_mask       : integer := 1;
        vc_alloc_type   : integer := 0;
        vc_alloc_arbiter_type: integer := 0;
        vc_alloc_prefer_empty: integer := 0;
        sw_alloc_type   : integer := 0;
        sw_alloc_arbiter_type: integer := 0;
        sw_alloc_spec_type: integer := 3;
        crossbar_type   : integer := 1;
        reset_type      : integer := 0;
        lfsr_index      : integer := 0;
        cfg_node_addr_width: integer := 10;
        cfg_reg_addr_width: integer := 6;
        cfg_data_width  : integer := 32;
        num_packets_width: integer := 16;
        arrival_rv_width: integer := 16;
        mc_idx_rv_width : integer := 4;
        rc_idx_rv_width : integer := 4;
        plength_idx_rv_width: integer := 4;
        num_plength_vals: integer := 2;
        packet_count_width: integer := 8;
        done_delay_width: integer := 6
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        io_node_addr_base: in     vl_logic_vector;
        io_write        : in     vl_logic;
        io_read         : in     vl_logic;
        io_addr         : in     vl_logic_vector;
        io_write_data   : in     vl_logic_vector;
        io_read_data    : out    vl_logic_vector;
        io_done         : out    vl_logic;
        error           : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of topology : constant is 1;
    attribute mti_svvh_generic_type of buffer_size : constant is 1;
    attribute mti_svvh_generic_type of num_message_classes : constant is 1;
    attribute mti_svvh_generic_type of num_resource_classes : constant is 1;
    attribute mti_svvh_generic_type of num_vcs_per_class : constant is 1;
    attribute mti_svvh_generic_type of num_nodes : constant is 1;
    attribute mti_svvh_generic_type of num_dimensions : constant is 1;
    attribute mti_svvh_generic_type of num_nodes_per_router : constant is 1;
    attribute mti_svvh_generic_type of packet_format : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_type : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_bypass : constant is 1;
    attribute mti_svvh_generic_type of max_payload_length : constant is 1;
    attribute mti_svvh_generic_type of min_payload_length : constant is 1;
    attribute mti_svvh_generic_type of router_type : constant is 1;
    attribute mti_svvh_generic_type of enable_link_pm : constant is 1;
    attribute mti_svvh_generic_type of flit_data_width : constant is 1;
    attribute mti_svvh_generic_type of error_capture_mode : constant is 1;
    attribute mti_svvh_generic_type of restrict_turns : constant is 1;
    attribute mti_svvh_generic_type of predecode_lar_info : constant is 1;
    attribute mti_svvh_generic_type of routing_type : constant is 1;
    attribute mti_svvh_generic_type of dim_order : constant is 1;
    attribute mti_svvh_generic_type of input_stage_can_hold : constant is 1;
    attribute mti_svvh_generic_type of fb_regfile_type : constant is 1;
    attribute mti_svvh_generic_type of fb_mgmt_type : constant is 1;
    attribute mti_svvh_generic_type of fb_fast_peek : constant is 1;
    attribute mti_svvh_generic_type of disable_static_reservations : constant is 1;
    attribute mti_svvh_generic_type of explicit_pipeline_register : constant is 1;
    attribute mti_svvh_generic_type of gate_buffer_write : constant is 1;
    attribute mti_svvh_generic_type of dual_path_alloc : constant is 1;
    attribute mti_svvh_generic_type of dual_path_allow_conflicts : constant is 1;
    attribute mti_svvh_generic_type of dual_path_mask_on_ready : constant is 1;
    attribute mti_svvh_generic_type of precomp_ivc_sel : constant is 1;
    attribute mti_svvh_generic_type of precomp_ip_sel : constant is 1;
    attribute mti_svvh_generic_type of elig_mask : constant is 1;
    attribute mti_svvh_generic_type of vc_alloc_type : constant is 1;
    attribute mti_svvh_generic_type of vc_alloc_arbiter_type : constant is 1;
    attribute mti_svvh_generic_type of vc_alloc_prefer_empty : constant is 1;
    attribute mti_svvh_generic_type of sw_alloc_type : constant is 1;
    attribute mti_svvh_generic_type of sw_alloc_arbiter_type : constant is 1;
    attribute mti_svvh_generic_type of sw_alloc_spec_type : constant is 1;
    attribute mti_svvh_generic_type of crossbar_type : constant is 1;
    attribute mti_svvh_generic_type of reset_type : constant is 1;
    attribute mti_svvh_generic_type of lfsr_index : constant is 1;
    attribute mti_svvh_generic_type of cfg_node_addr_width : constant is 1;
    attribute mti_svvh_generic_type of cfg_reg_addr_width : constant is 1;
    attribute mti_svvh_generic_type of cfg_data_width : constant is 1;
    attribute mti_svvh_generic_type of num_packets_width : constant is 1;
    attribute mti_svvh_generic_type of arrival_rv_width : constant is 1;
    attribute mti_svvh_generic_type of mc_idx_rv_width : constant is 1;
    attribute mti_svvh_generic_type of rc_idx_rv_width : constant is 1;
    attribute mti_svvh_generic_type of plength_idx_rv_width : constant is 1;
    attribute mti_svvh_generic_type of num_plength_vals : constant is 1;
    attribute mti_svvh_generic_type of packet_count_width : constant is 1;
    attribute mti_svvh_generic_type of done_delay_width : constant is 1;
end tc_router_wrap;
