library verilog;
use verilog.vl_types.all;
entity whr_ip_ctrl_mac is
    generic(
        buffer_size     : integer := 8;
        num_routers_per_dim: integer := 4;
        num_dimensions  : integer := 2;
        num_nodes_per_router: integer := 1;
        connectivity    : integer := 0;
        packet_format   : integer := 2;
        flow_ctrl_type  : integer := 0;
        elig_mask       : integer := 0;
        max_payload_length: integer := 4;
        min_payload_length: integer := 1;
        enable_link_pm  : integer := 1;
        flit_data_width : integer := 64;
        restrict_turns  : integer := 1;
        routing_type    : integer := 0;
        dim_order       : integer := 0;
        input_stage_can_hold: integer := 0;
        fb_regfile_type : integer := 0;
        fb_fast_peek    : integer := 1;
        explicit_pipeline_register: integer := 0;
        gate_buffer_write: integer := 0;
        error_capture_mode: integer := 1;
        port_id         : integer := 0;
        reset_type      : integer := 0
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        router_address  : in     vl_logic_vector;
        channel_in      : in     vl_logic_vector;
        route_op        : out    vl_logic_vector;
        req             : out    vl_logic;
        req_head        : out    vl_logic;
        req_tail        : out    vl_logic;
        gnt             : in     vl_logic;
        flit_data_out   : out    vl_logic_vector;
        flow_ctrl_out   : out    vl_logic_vector;
        error           : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of buffer_size : constant is 1;
    attribute mti_svvh_generic_type of num_routers_per_dim : constant is 1;
    attribute mti_svvh_generic_type of num_dimensions : constant is 1;
    attribute mti_svvh_generic_type of num_nodes_per_router : constant is 1;
    attribute mti_svvh_generic_type of connectivity : constant is 1;
    attribute mti_svvh_generic_type of packet_format : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_type : constant is 1;
    attribute mti_svvh_generic_type of elig_mask : constant is 1;
    attribute mti_svvh_generic_type of max_payload_length : constant is 1;
    attribute mti_svvh_generic_type of min_payload_length : constant is 1;
    attribute mti_svvh_generic_type of enable_link_pm : constant is 1;
    attribute mti_svvh_generic_type of flit_data_width : constant is 1;
    attribute mti_svvh_generic_type of restrict_turns : constant is 1;
    attribute mti_svvh_generic_type of routing_type : constant is 1;
    attribute mti_svvh_generic_type of dim_order : constant is 1;
    attribute mti_svvh_generic_type of input_stage_can_hold : constant is 1;
    attribute mti_svvh_generic_type of fb_regfile_type : constant is 1;
    attribute mti_svvh_generic_type of fb_fast_peek : constant is 1;
    attribute mti_svvh_generic_type of explicit_pipeline_register : constant is 1;
    attribute mti_svvh_generic_type of gate_buffer_write : constant is 1;
    attribute mti_svvh_generic_type of error_capture_mode : constant is 1;
    attribute mti_svvh_generic_type of port_id : constant is 1;
    attribute mti_svvh_generic_type of reset_type : constant is 1;
end whr_ip_ctrl_mac;
