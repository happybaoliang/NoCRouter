library verilog;
use verilog.vl_types.all;
entity rtr_alloc_mac is
    generic(
        num_message_classes: integer := 2;
        num_resource_classes: integer := 2;
        num_vcs_per_class: integer := 1;
        num_routers_per_dim: integer := 4;
        num_dimensions  : integer := 2;
        num_nodes_per_router: integer := 1;
        connectivity    : integer := 0;
        flow_ctrl_type  : integer := 0;
        restrict_turns  : integer := 1;
        routing_type    : integer := 0;
        dim_order       : integer := 0;
        precomp_ivc_sel : integer := 1;
        precomp_ip_sel  : integer := 1;
        fb_mgmt_type    : integer := 0;
        elig_mask       : integer := 0;
        sw_alloc_arbiter_type: integer := 0;
        vc_alloc_arbiter_type: integer := 0;
        vc_alloc_prefer_empty: integer := 0;
        dual_path_alloc : integer := 1;
        dual_path_allow_conflicts: integer := 0;
        dual_path_mask_on_ready: integer := 1;
        reset_type      : integer := 0
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        route_in_ip_ivc_op: in     vl_logic_vector;
        route_in_ip_ivc_orc: in     vl_logic_vector;
        flit_valid_in_ip_ivc: in     vl_logic_vector;
        flit_last_in_ip_ivc: in     vl_logic_vector;
        flit_head_in_ip_ivc: in     vl_logic_vector;
        flit_tail_in_ip_ivc: in     vl_logic_vector;
        route_fast_in_ip_op: in     vl_logic_vector;
        route_fast_in_ip_orc: in     vl_logic_vector;
        flit_valid_fast_in_ip: in     vl_logic_vector;
        flit_head_fast_in_ip: in     vl_logic_vector;
        flit_tail_fast_in_ip: in     vl_logic_vector;
        flit_sel_fast_in_ip_ivc: in     vl_logic_vector;
        flit_sel_out_ip_ivc: out    vl_logic_vector;
        flit_sent_out_ip: out    vl_logic_vector;
        flit_sel_fast_out_ip: out    vl_logic_vector;
        flit_sent_fast_out_ip: out    vl_logic_vector;
        flit_sel_out_op_ip: out    vl_logic_vector;
        flit_valid_out_op: out    vl_logic_vector;
        flit_head_out_op: out    vl_logic_vector;
        flit_tail_out_op: out    vl_logic_vector;
        flit_sel_out_op_ovc: out    vl_logic_vector;
        elig_in_op_ovc  : in     vl_logic_vector;
        empty_in_op_ovc : in     vl_logic_vector;
        almost_full_in_op_ovc: in     vl_logic_vector;
        full_in_op_ovc  : in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of num_message_classes : constant is 1;
    attribute mti_svvh_generic_type of num_resource_classes : constant is 1;
    attribute mti_svvh_generic_type of num_vcs_per_class : constant is 1;
    attribute mti_svvh_generic_type of num_routers_per_dim : constant is 1;
    attribute mti_svvh_generic_type of num_dimensions : constant is 1;
    attribute mti_svvh_generic_type of num_nodes_per_router : constant is 1;
    attribute mti_svvh_generic_type of connectivity : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_type : constant is 1;
    attribute mti_svvh_generic_type of restrict_turns : constant is 1;
    attribute mti_svvh_generic_type of routing_type : constant is 1;
    attribute mti_svvh_generic_type of dim_order : constant is 1;
    attribute mti_svvh_generic_type of precomp_ivc_sel : constant is 1;
    attribute mti_svvh_generic_type of precomp_ip_sel : constant is 1;
    attribute mti_svvh_generic_type of fb_mgmt_type : constant is 1;
    attribute mti_svvh_generic_type of elig_mask : constant is 1;
    attribute mti_svvh_generic_type of sw_alloc_arbiter_type : constant is 1;
    attribute mti_svvh_generic_type of vc_alloc_arbiter_type : constant is 1;
    attribute mti_svvh_generic_type of vc_alloc_prefer_empty : constant is 1;
    attribute mti_svvh_generic_type of dual_path_alloc : constant is 1;
    attribute mti_svvh_generic_type of dual_path_allow_conflicts : constant is 1;
    attribute mti_svvh_generic_type of dual_path_mask_on_ready : constant is 1;
    attribute mti_svvh_generic_type of reset_type : constant is 1;
end rtr_alloc_mac;
