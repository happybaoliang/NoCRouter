library verilog;
use verilog.vl_types.all;
entity vcr_ivc_ctrl is
    generic(
        num_message_classes: integer := 2;
        num_resource_classes: integer := 2;
        num_vcs_per_class: integer := 1;
        num_routers_per_dim: integer := 4;
        num_dimensions  : integer := 2;
        num_nodes_per_router: integer := 1;
        connectivity    : integer := 0;
        packet_format   : integer := 2;
        max_payload_length: integer := 4;
        min_payload_length: integer := 1;
        restrict_turns  : integer := 1;
        routing_type    : integer := 0;
        dim_order       : integer := 0;
        elig_mask       : integer := 0;
        sw_alloc_spec   : integer := 1;
        fb_mgmt_type    : integer := 0;
        explicit_pipeline_register: integer := 0;
        vc_id           : integer := 0;
        port_id         : integer := 0;
        reset_type      : integer := 0
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        router_address  : in     vl_logic_vector;
        flit_valid_in   : in     vl_logic;
        flit_head_in    : in     vl_logic;
        flit_tail_in    : in     vl_logic;
        flit_sel_in     : in     vl_logic;
        header_info_in  : in     vl_logic_vector;
        fb_pop_tail     : in     vl_logic;
        fb_pop_next_header_info: in     vl_logic_vector;
        almost_full_op_ovc: in     vl_logic_vector;
        full_op_ovc     : in     vl_logic_vector;
        route_op        : out    vl_logic_vector;
        route_orc       : out    vl_logic_vector;
        vc_gnt          : in     vl_logic;
        vc_sel_ovc      : in     vl_logic_vector;
        sw_gnt          : in     vl_logic;
        sw_sel          : in     vl_logic;
        sw_gnt_op       : in     vl_logic_vector;
        flit_valid      : out    vl_logic;
        flit_head       : out    vl_logic;
        flit_tail       : out    vl_logic;
        next_lar_info   : out    vl_logic_vector;
        fb_almost_empty : in     vl_logic;
        fb_empty        : in     vl_logic;
        allocated       : out    vl_logic;
        free_nonspec    : out    vl_logic;
        free_spec       : out    vl_logic;
        errors          : out    vl_logic_vector(0 to 2)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of num_message_classes : constant is 1;
    attribute mti_svvh_generic_type of num_resource_classes : constant is 1;
    attribute mti_svvh_generic_type of num_vcs_per_class : constant is 1;
    attribute mti_svvh_generic_type of num_routers_per_dim : constant is 1;
    attribute mti_svvh_generic_type of num_dimensions : constant is 1;
    attribute mti_svvh_generic_type of num_nodes_per_router : constant is 1;
    attribute mti_svvh_generic_type of connectivity : constant is 1;
    attribute mti_svvh_generic_type of packet_format : constant is 1;
    attribute mti_svvh_generic_type of max_payload_length : constant is 1;
    attribute mti_svvh_generic_type of min_payload_length : constant is 1;
    attribute mti_svvh_generic_type of restrict_turns : constant is 1;
    attribute mti_svvh_generic_type of routing_type : constant is 1;
    attribute mti_svvh_generic_type of dim_order : constant is 1;
    attribute mti_svvh_generic_type of elig_mask : constant is 1;
    attribute mti_svvh_generic_type of sw_alloc_spec : constant is 1;
    attribute mti_svvh_generic_type of fb_mgmt_type : constant is 1;
    attribute mti_svvh_generic_type of explicit_pipeline_register : constant is 1;
    attribute mti_svvh_generic_type of vc_id : constant is 1;
    attribute mti_svvh_generic_type of port_id : constant is 1;
    attribute mti_svvh_generic_type of reset_type : constant is 1;
end vcr_ivc_ctrl;
