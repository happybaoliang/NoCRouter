library verilog;
use verilog.vl_types.all;
entity rtr_top is
    generic(
        buffer_size     : integer := 32;
        num_message_classes: integer := 2;
        num_resource_classes: integer := 2;
        num_vcs_per_class: integer := 1;
        num_routers_per_dim: integer := 4;
        num_dimensions  : integer := 2;
        num_nodes_per_router: integer := 1;
        connectivity    : integer := 0;
        packet_format   : integer := 2;
        flow_ctrl_type  : integer := 0;
        flow_ctrl_bypass: integer := 1;
        max_payload_length: integer := 4;
        min_payload_length: integer := 1;
        enable_link_pm  : integer := 1;
        flit_data_width : integer := 64;
        error_capture_mode: integer := 1;
        restrict_turns  : integer := 1;
        predecode_lar_info: integer := 1;
        routing_type    : integer := 0;
        dim_order       : integer := 0;
        fb_regfile_type : integer := 0;
        fb_mgmt_type    : integer := 0;
        fb_fast_peek    : integer := 1;
        disable_static_reservations: integer := 0;
        explicit_pipeline_register: integer := 0;
        gate_buffer_write: integer := 0;
        dual_path_alloc : integer := 1;
        dual_path_allow_conflicts: integer := 0;
        dual_path_mask_on_ready: integer := 1;
        precomp_ivc_sel : integer := 1;
        precomp_ip_sel  : integer := 1;
        elig_mask       : integer := 0;
        sw_alloc_arbiter_type: integer := 0;
        vc_alloc_arbiter_type: integer := 0;
        vc_alloc_prefer_empty: integer := 0;
        crossbar_type   : integer := 1;
        reset_type      : integer := 0
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        router_address  : in     vl_logic_vector;
        channel_in_ip   : in     vl_logic_vector;
        flow_ctrl_out_ip: out    vl_logic_vector;
        channel_out_op  : out    vl_logic_vector;
        flow_ctrl_in_op : in     vl_logic_vector;
        error           : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of buffer_size : constant is 1;
    attribute mti_svvh_generic_type of num_message_classes : constant is 1;
    attribute mti_svvh_generic_type of num_resource_classes : constant is 1;
    attribute mti_svvh_generic_type of num_vcs_per_class : constant is 1;
    attribute mti_svvh_generic_type of num_routers_per_dim : constant is 1;
    attribute mti_svvh_generic_type of num_dimensions : constant is 1;
    attribute mti_svvh_generic_type of num_nodes_per_router : constant is 1;
    attribute mti_svvh_generic_type of connectivity : constant is 1;
    attribute mti_svvh_generic_type of packet_format : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_type : constant is 1;
    attribute mti_svvh_generic_type of flow_ctrl_bypass : constant is 1;
    attribute mti_svvh_generic_type of max_payload_length : constant is 1;
    attribute mti_svvh_generic_type of min_payload_length : constant is 1;
    attribute mti_svvh_generic_type of enable_link_pm : constant is 1;
    attribute mti_svvh_generic_type of flit_data_width : constant is 1;
    attribute mti_svvh_generic_type of error_capture_mode : constant is 1;
    attribute mti_svvh_generic_type of restrict_turns : constant is 1;
    attribute mti_svvh_generic_type of predecode_lar_info : constant is 1;
    attribute mti_svvh_generic_type of routing_type : constant is 1;
    attribute mti_svvh_generic_type of dim_order : constant is 1;
    attribute mti_svvh_generic_type of fb_regfile_type : constant is 1;
    attribute mti_svvh_generic_type of fb_mgmt_type : constant is 1;
    attribute mti_svvh_generic_type of fb_fast_peek : constant is 1;
    attribute mti_svvh_generic_type of disable_static_reservations : constant is 1;
    attribute mti_svvh_generic_type of explicit_pipeline_register : constant is 1;
    attribute mti_svvh_generic_type of gate_buffer_write : constant is 1;
    attribute mti_svvh_generic_type of dual_path_alloc : constant is 1;
    attribute mti_svvh_generic_type of dual_path_allow_conflicts : constant is 1;
    attribute mti_svvh_generic_type of dual_path_mask_on_ready : constant is 1;
    attribute mti_svvh_generic_type of precomp_ivc_sel : constant is 1;
    attribute mti_svvh_generic_type of precomp_ip_sel : constant is 1;
    attribute mti_svvh_generic_type of elig_mask : constant is 1;
    attribute mti_svvh_generic_type of sw_alloc_arbiter_type : constant is 1;
    attribute mti_svvh_generic_type of vc_alloc_arbiter_type : constant is 1;
    attribute mti_svvh_generic_type of vc_alloc_prefer_empty : constant is 1;
    attribute mti_svvh_generic_type of crossbar_type : constant is 1;
    attribute mti_svvh_generic_type of reset_type : constant is 1;
end rtr_top;
